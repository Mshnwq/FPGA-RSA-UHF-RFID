module dataPath
	#(parameter WordSize = 8)
	(  
	input clk, reset,
	
	// Data Path I/O	
	input  [WordSize-1:0] input_text,
	input  [WordSize-1:0] key,
	output [WordSize-1:0] output_text,
	
	// Controller I/O
	input wire go,       // enablers
	output wire done     // flags
	);
	

endmodule 